module GameBoard   ( input              clk, reset
                     input logic [11:0] piecesIn [64],
						   output logic [11:0] piecesOut [64]);
							
	always_ff @ (posedge clk)
    case (reset)
		1'b1: begin 
			piecesOut <= {12'b000000000100, 12'b000000010000, 12'b000000001000, 12'b000000000010, 12'b000000000001, 12'b000000001000, 12'b000000010000, 12'b000000000100,
							  12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000,
							  12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000,
							  12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000,
							  12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000,
							  12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000,
							  12'b100000000000, 12'b100000000000, 12'b100000000000, 12'b100000000000, 12'b100000000000, 12'b100000000000, 12'b100000000000, 12'b100000000000,
							  12'b000100000000, 12'b010000000000, 12'b001000000000, 12'b000010000000, 12'b000001000000, 12'b001000000000, 12'b010000000000, 12'b000100000000} 
		end    
		default: begin
			piecesOut <= piecesIn;
		end 
	 
    endcase						
endmodule 